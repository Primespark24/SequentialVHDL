-----------------------------------------------
-- Module Name:    divideby3FSM 
-- A true divide by 3 clock with 50% duty cycle
-----------------------------------------------
library IEEE; use IEEE.STD_LOGIC_1164.ALL;

entity divideby3FSM_50 is
    port ( clk :   in  STD_LOGIC;
           reset : in  STD_LOGIC;
           y :    out  STD_LOGIC);
end divideby3FSM_50;

architecture Behavioral of divideby3FSM_50 is
	-- create signals here to wire the hardware edge
	-- triggered latches together
begin

   -- Edge Triggered Latch A goes here

   -- Edge Triggered Latch B goes here
	
   -- Edge Triggered Latch C goes here

   -- Generate the output signal y here
	
end Behavioral;